library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package wave_rom_package is
	type wave_rom_logic_vector_array is array (1023 downto 0) of std_logic_vector (31 downto 0);
	type wave_rom_unsigned_array is array (1023 downto 0) of Unsigned (31 downto 0);

	signal rom_core: wave_rom_logic_vector_array:=(
		0	 => "00000000000000000000000000000000",
		1	 => "00000000001100100100001111110101",
		2	 => "00000000011001001000011111100010",
		3	 => "00000000100101101100101111000001",
		4	 => "00000000110010010000111110000111",
		5	 => "00000000111110110101001100101111",
		6	 => "00000001001011011001011010110000",
		7	 => "00000001010111111101101000000011",
		8	 => "00000001100100100001110100011111",
		9	 => "00000001110001000101111111111110",
		10	 => "00000001111101101010001010010110",
		11	 => "00000010001010001110010011100001",
		12	 => "00000010010110110010011011010111",
		13	 => "00000010100011010110100001110000",
		14	 => "00000010101111111010100110100100",
		15	 => "00000010111100011110101001101011",
		16	 => "00000011001001000010101010111110",
		17	 => "00000011010101100110101010010110",
		18	 => "00000011100010001010100111101001",
		19	 => "00000011101110101110100010110001",
		20	 => "00000011111011010010011011100110",
		21	 => "00000100000111110110010001111111",
		22	 => "00000100010100011010000101110110",
		23	 => "00000100100000111101110111000011",
		24	 => "00000100101101100001100101011101",
		25	 => "00000100111010000101010000111101",
		26	 => "00000101000110101000111001011011",
		27	 => "00000101010011001100011110110000",
		28	 => "00000101011111110000000000110100",
		29	 => "00000101101100010011011111011111",
		30	 => "00000101111000110110111010101001",
		31	 => "00000110000101011010010010001010",
		32	 => "00000110010001111101100101111100",
		33	 => "00000110011110100000110101110101",
		34	 => "00000110101011000100000001101111",
		35	 => "00000110110111100111001001100001",
		36	 => "00000111000100001010001101000100",
		37	 => "00000111010000101101001100010000",
		38	 => "00000111011101010000000110111110",
		39	 => "00000111101001110010111101000101",
		40	 => "00000111110110010101101110011110",
		41	 => "00001000000010111000011011000001",
		42	 => "00001000001111011011000010100111",
		43	 => "00001000011011111101100101000111",
		44	 => "00001000101000100000000010011010",
		45	 => "00001000110101000010011010011000",
		46	 => "00001001000001100100101100111010",
		47	 => "00001001001110000110111001110111",
		48	 => "00001001011010101001000001001001",
		49	 => "00001001100111001011000010100111",
		50	 => "00001001110011101100111110001001",
		51	 => "00001010000000001110110011101000",
		52	 => "00001010001100110000100010111100",
		53	 => "00001010011001010010001011111110",
		54	 => "00001010100101110011101110100101",
		55	 => "00001010110010010101001010101010",
		56	 => "00001010111110110110100000000101",
		57	 => "00001011001011010111101110101110",
		58	 => "00001011010111111000110110011111",
		59	 => "00001011100100011001110111001110",
		60	 => "00001011110000111010110000110101",
		61	 => "00001011111101011011100011001011",
		62	 => "00001100001001111100001110001001",
		63	 => "00001100010110011100110001100111",
		64	 => "00001100100010111101001101011110",
		65	 => "00001100101111011101100001100101",
		66	 => "00001100111011111101101101110101",
		67	 => "00001101001000011101110010000111",
		68	 => "00001101010100111101101110010010",
		69	 => "00001101100001011101100010001111",
		70	 => "00001101101101111101001101110110",
		71	 => "00001101111010011100110000111111",
		72	 => "00001110000110111100001011100011",
		73	 => "00001110010011011011011101011011",
		74	 => "00001110011111111010100110011101",
		75	 => "00001110101100011001100110100011",
		76	 => "00001110111000111000011101100101",
		77	 => "00001111000101010111001011011100",
		78	 => "00001111010001110101101111111110",
		79	 => "00001111011110010100001011000110",
		80	 => "00001111101010110010011100101011",
		81	 => "00001111110111010000100100100101",
		82	 => "00010000000011101110100010101101",
		83	 => "00010000010000001100010110111011",
		84	 => "00010000011100101010000001000111",
		85	 => "00010000101001000111100001001010",
		86	 => "00010000110101100100110110111100",
		87	 => "00010001000010000010000010010101",
		88	 => "00010001001110011111000011001110",
		89	 => "00010001011010111011111001011111",
		90	 => "00010001100111011000100101000000",
		91	 => "00010001110011110101000101101010",
		92	 => "00010010000000010001011011010100",
		93	 => "00010010001100101101100101111000",
		94	 => "00010010011001001001100101001101",
		95	 => "00010010100101100101011001001101",
		96	 => "00010010110010000001000001101110",
		97	 => "00010010111110011100011110101010",
		98	 => "00010011001010110111101111111001",
		99	 => "00010011010111010010110101010011",
		100	 => "00010011100011101101101110110000",
		101	 => "00010011110000001000011100001010",
		102	 => "00010011111100100010111101010111",
		103	 => "00010100001000111101010010010010",
		104	 => "00010100010101010111011010110001",
		105	 => "00010100100001110001010110101101",
		106	 => "00010100101110001011000101111111",
		107	 => "00010100111010100100101000011111",
		108	 => "00010101000110111101111110000101",
		109	 => "00010101010011010111000110101010",
		110	 => "00010101011111110000000010000110",
		111	 => "00010101101100001000110000010001",
		112	 => "00010101111000100001010001000100",
		113	 => "00010110000100111001100100010111",
		114	 => "00010110010001010001101010000011",
		115	 => "00010110011101101001100001111111",
		116	 => "00010110101010000001001100000100",
		117	 => "00010110110110011000101000001100",
		118	 => "00010111000010101111110110001101",
		119	 => "00010111001111000110110110000000",
		120	 => "00010111011011011101100111011110",
		121	 => "00010111100111110100001010011111",
		122	 => "00010111110100001010011110111011",
		123	 => "00011000000000100000100100101100",
		124	 => "00011000001100110110011011101000",
		125	 => "00011000011001001100000011101001",
		126	 => "00011000100101100001011100100111",
		127	 => "00011000110001110110100110011011",
		128	 => "00011000111110001011100000111100",
		129	 => "00011001001010100000001100000011",
		130	 => "00011001010110110100100111101001",
		131	 => "00011001100011001000110011100110",
		132	 => "00011001101111011100101111110010",
		133	 => "00011001111011110000011100000110",
		134	 => "00011010001000000011111000011011",
		135	 => "00011010010100010111000100100111",
		136	 => "00011010100000101010000000100101",
		137	 => "00011010101100111100101100001100",
		138	 => "00011010111001001111000111010101",
		139	 => "00011011000101100001010001111001",
		140	 => "00011011010001110011001011101111",
		141	 => "00011011011110000100110100110000",
		142	 => "00011011101010010110001100110100",
		143	 => "00011011110110100111010011110101",
		144	 => "00011100000010111000001001101010",
		145	 => "00011100001111001000101110001100",
		146	 => "00011100011011011001000001010011",
		147	 => "00011100100111101001000010111000",
		148	 => "00011100110011111000110010110011",
		149	 => "00011101000000001000010000111100",
		150	 => "00011101001100010111011101001101",
		151	 => "00011101011000100110010111011101",
		152	 => "00011101100100110100111111100101",
		153	 => "00011101110001000011010101011101",
		154	 => "00011101111101010001011000111111",
		155	 => "00011110001001011111001010000001",
		156	 => "00011110010101101100101000011110",
		157	 => "00011110100001111001110100001100",
		158	 => "00011110101110000110101101000110",
		159	 => "00011110111010010011010011000010",
		160	 => "00011111000110011111100101111011",
		161	 => "00011111010010101011100101100111",
		162	 => "00011111011110110111010010000000",
		163	 => "00011111101011000010101010111110",
		164	 => "00011111110111001101110000011010",
		165	 => "00100000000011011000100010001100",
		166	 => "00100000001111100011000000001101",
		167	 => "00100000011011101101001010010101",
		168	 => "00100000100111110111000000011100",
		169	 => "00100000110100000000100010011011",
		170	 => "00100001000000001001110000001011",
		171	 => "00100001001100010010101001100100",
		172	 => "00100001011000011011001110011111",
		173	 => "00100001100100100011011110110100",
		174	 => "00100001110000101011011010011100",
		175	 => "00100001111100110011000001001110",
		176	 => "00100010001000111010010011000101",
		177	 => "00100010010101000001001111111000",
		178	 => "00100010100001000111110111011111",
		179	 => "00100010101101001110001001110100",
		180	 => "00100010111001010100000110101110",
		181	 => "00100011000101011001101110000111",
		182	 => "00100011010001011110111111110111",
		183	 => "00100011011101100011111011110111",
		184	 => "00100011101001101000100001111110",
		185	 => "00100011110101101100110010000110",
		186	 => "00100100000001110000101100000111",
		187	 => "00100100001101110100001111111010",
		188	 => "00100100011001110111011101010111",
		189	 => "00100100100101111010010100010111",
		190	 => "00100100110001111100110100110010",
		191	 => "00100100111101111110111110100001",
		192	 => "00100101001010000000110001011101",
		193	 => "00100101010110000010001101011110",
		194	 => "00100101100010000011010010011101",
		195	 => "00100101101110000100000000010010",
		196	 => "00100101111010000100010110110101",
		197	 => "00100110000110000100010110000001",
		198	 => "00100110010010000011111101101100",
		199	 => "00100110011110000011001101110000",
		200	 => "00100110101010000010000110000101",
		201	 => "00100110110110000000100110100100",
		202	 => "00100111000001111110101111000110",
		203	 => "00100111001101111100011111100011",
		204	 => "00100111011001111001110111110100",
		205	 => "00100111100101110110110111110000",
		206	 => "00100111110001110011011111010010",
		207	 => "00100111111101101111101110010010",
		208	 => "00101000001001101011100100101000",
		209	 => "00101000010101100111000010001100",
		210	 => "00101000100001100010000110111001",
		211	 => "00101000101101011100110010100101",
		212	 => "00101000111001010111000101001010",
		213	 => "00101001000101010000111110100001",
		214	 => "00101001010001001010011110100010",
		215	 => "00101001011101000011100101000101",
		216	 => "00101001101000111100010010000100",
		217	 => "00101001110100110100100101011000",
		218	 => "00101010000000101100011110111000",
		219	 => "00101010001100100011111110011101",
		220	 => "00101010011000011011000100000001",
		221	 => "00101010100100010001101111011011",
		222	 => "00101010110000001000000000100101",
		223	 => "00101010111011111101110111011000",
		224	 => "00101011000111110011010011101011",
		225	 => "00101011010011101000010101011000",
		226	 => "00101011011111011100111100010111",
		227	 => "00101011101011010001001000100001",
		228	 => "00101011110111000100111001101111",
		229	 => "00101100000010111000001111111001",
		230	 => "00101100001110101011001010111001",
		231	 => "00101100011010011101101010100110",
		232	 => "00101100100110001111101110111010",
		233	 => "00101100110010000001010111101101",
		234	 => "00101100111101110010100100111001",
		235	 => "00101101001001100011010110010101",
		236	 => "00101101010101010011101011111011",
		237	 => "00101101100001000011100101100011",
		238	 => "00101101101100110011000011000111",
		239	 => "00101101111000100010000100011110",
		240	 => "00101110000100010000101001100001",
		241	 => "00101110001111111110110010001011",
		242	 => "00101110011011101100011110010010",
		243	 => "00101110100111011001101101110000",
		244	 => "00101110110011000110100000011110",
		245	 => "00101110111110110010110110010100",
		246	 => "00101111001010011110101111001100",
		247	 => "00101111010110001010001010111101",
		248	 => "00101111100001110101001001100010",
		249	 => "00101111101101011111101010110010",
		250	 => "00101111111001001001101110100110",
		251	 => "00110000000100110011010100111000",
		252	 => "00110000010000011100011101100000",
		253	 => "00110000011100000101001000010111",
		254	 => "00110000100111101101010101010101",
		255	 => "00110000110011010101000100010100",
		256	 => "00110000111110111100010101001101",
		257	 => "00110001001010100011000111110111",
		258	 => "00110001010110001001011100001101",
		259	 => "00110001100001101111010010000111",
		260	 => "00110001101101010100101001011101",
		261	 => "00110001111000111001100010001001",
		262	 => "00110010000100011101111100000011",
		263	 => "00110010010000000001110111000101",
		264	 => "00110010011011100101010011000111",
		265	 => "00110010100111001000010000000010",
		266	 => "00110010110010101010101101101111",
		267	 => "00110010111110001100101100000111",
		268	 => "00110011001001101110001011000010",
		269	 => "00110011010101001111001010011010",
		270	 => "00110011100000101111101010001000",
		271	 => "00110011101100001111101010000100",
		272	 => "00110011110111101111001010000111",
		273	 => "00110100000011001110001010001010",
		274	 => "00110100001110101100101010000111",
		275	 => "00110100011010001010101001110110",
		276	 => "00110100100101101000001001001111",
		277	 => "00110100110001000101001000001101",
		278	 => "00110100111100100001100110100111",
		279	 => "00110101000111111101100100010111",
		280	 => "00110101010011011001000001010110",
		281	 => "00110101011110110011111101011101",
		282	 => "00110101101010001110011000100100",
		283	 => "00110101110101101000010010100101",
		284	 => "00110110000001000001101011011000",
		285	 => "00110110001100011010100010110111",
		286	 => "00110110010111110010111000111011",
		287	 => "00110110100011001010101101011100",
		288	 => "00110110101110100010000000010011",
		289	 => "00110110111001111000110001011010",
		290	 => "00110111000101001111000000101001",
		291	 => "00110111010000100100101101111010",
		292	 => "00110111011011111001111001000110",
		293	 => "00110111100111001110100010000100",
		294	 => "00110111110010100010101000101111",
		295	 => "00110111111101110110001101000000",
		296	 => "00111000001001001001001110110000",
		297	 => "00111000010100011011101101110110",
		298	 => "00111000011111101101101010001110",
		299	 => "00111000101010111111000011101111",
		300	 => "00111000110110001111111010010011",
		301	 => "00111001000001100000001101110010",
		302	 => "00111001001100101111111110000111",
		303	 => "00111001010111111111001011001001",
		304	 => "00111001100011001101110100110010",
		305	 => "00111001101110011011111010111011",
		306	 => "00111001111001101001011101011101",
		307	 => "00111010000100110110011100010010",
		308	 => "00111010010000000010110111010001",
		309	 => "00111010011011001110101110010101",
		310	 => "00111010100110011010000001010111",
		311	 => "00111010110001100100110000001111",
		312	 => "00111010111100101110111010110111",
		313	 => "00111011000111111000100001000111",
		314	 => "00111011010011000001100010111001",
		315	 => "00111011011110001010000000000111",
		316	 => "00111011101001010001111000101001",
		317	 => "00111011110100011001001100010111",
		318	 => "00111011111111011111111011001101",
		319	 => "00111100001010100110000101000010",
		320	 => "00111100010101101011101001110000",
		321	 => "00111100100000110000101001001111",
		322	 => "00111100101011110101000011011010",
		323	 => "00111100110110111000111000001001",
		324	 => "00111101000001111100000111010101",
		325	 => "00111101001100111110110000111001",
		326	 => "00111101011000000000110100101011",
		327	 => "00111101100011000010010010100111",
		328	 => "00111101101110000011001010100101",
		329	 => "00111101111001000011011100011111",
		330	 => "00111110000100000011001000001101",
		331	 => "00111110001111000010001101101001",
		332	 => "00111110011010000000101100101100",
		333	 => "00111110100100111110100101001111",
		334	 => "00111110101111111011110111001100",
		335	 => "00111110111010111000100010011100",
		336	 => "00111111000101110100100110110111",
		337	 => "00111111010000110000000100011000",
		338	 => "00111111011011101010111010111000",
		339	 => "00111111100110100101001010001111",
		340	 => "00111111110001011110110010010111",
		341	 => "00111111111100010111110011001010",
		342	 => "01000000000111010000001100100000",
		343	 => "01000000010010000111111110010011",
		344	 => "01000000011100111111001000011101",
		345	 => "01000000100111110101101010110110",
		346	 => "01000000110010101011100101010111",
		347	 => "01000000111101100000110111111011",
		348	 => "01000001001000010101100010011010",
		349	 => "01000001010011001001100100101110",
		350	 => "01000001011101111100111110110000",
		351	 => "01000001101000101111110000011010",
		352	 => "01000001110011100001111001100100",
		353	 => "01000001111110010011011010001000",
		354	 => "01000010001001000100010010000000",
		355	 => "01000010010011110100100001000101",
		356	 => "01000010011110100100000111010000",
		357	 => "01000010101001010011000100011010",
		358	 => "01000010110100000001011000011110",
		359	 => "01000010111110101111000011010011",
		360	 => "01000011001001011100000100110101",
		361	 => "01000011010100001000011100111100",
		362	 => "01000011011110110100001011100001",
		363	 => "01000011101001011111010000011110",
		364	 => "01000011110100001001101011101100",
		365	 => "01000011111110110011011101000101",
		366	 => "01000100001001011100100100100011",
		367	 => "01000100010100000101000001111110",
		368	 => "01000100011110101100110101010000",
		369	 => "01000100101001010011111110010011",
		370	 => "01000100110011111010011100111111",
		371	 => "01000100111110100000010001001111",
		372	 => "01000101001001000101011010111100",
		373	 => "01000101010011101001111010000000",
		374	 => "01000101011110001101101110010011",
		375	 => "01000101101000110000110111110000",
		376	 => "01000101110011010011010110001111",
		377	 => "01000101111101110101001001101011",
		378	 => "01000110001000010110010001111100",
		379	 => "01000110010010110110101110111101",
		380	 => "01000110011101010110100000100111",
		381	 => "01000110100111110101100110110100",
		382	 => "01000110110010010100000001011100",
		383	 => "01000110111100110001110000011010",
		384	 => "01000111000111001110110011100110",
		385	 => "01000111010001101011001010111100",
		386	 => "01000111011100000110110110010011",
		387	 => "01000111100110100001110101100110",
		388	 => "01000111110000111100001000101110",
		389	 => "01000111111011010101101111100110",
		390	 => "01001000000101101110101010000101",
		391	 => "01001000010000000110111000000111",
		392	 => "01001000011010011110011001100100",
		393	 => "01001000100100110101001110010111",
		394	 => "01001000101111001011010110011000",
		395	 => "01001000111001100000110001100010",
		396	 => "01001001000011110101011111101110",
		397	 => "01001001001110001001100000110101",
		398	 => "01001001011000011100110100110010",
		399	 => "01001001100010101111011011011110",
		400	 => "01001001101101000001010100110011",
		401	 => "01001001110111010010100000101010",
		402	 => "01001010000001100010111110111101",
		403	 => "01001010001011110010101111100101",
		404	 => "01001010010110000001110010011101",
		405	 => "01001010100000010000000111011110",
		406	 => "01001010101010011101101110100001",
		407	 => "01001010110100101010100111100001",
		408	 => "01001010111110110110110010010111",
		409	 => "01001011001001000010001110111101",
		410	 => "01001011010011001100111101001101",
		411	 => "01001011011101010110111100111111",
		412	 => "01001011100111100000001110001111",
		413	 => "01001011110001101000110000110110",
		414	 => "01001011111011110000100100101101",
		415	 => "01001100000101110111101001101110",
		416	 => "01001100001111111101111111110011",
		417	 => "01001100011010000011100110110110",
		418	 => "01001100100100001000011110110001",
		419	 => "01001100101110001100100111011101",
		420	 => "01001100111000010000000000110100",
		421	 => "01001101000010010010101010110000",
		422	 => "01001101001100010100100101001011",
		423	 => "01001101010110010101101111111110",
		424	 => "01001101100000010110001011000100",
		425	 => "01001101101010010101110110010110",
		426	 => "01001101110100010100110001101110",
		427	 => "01001101111110010010111101000101",
		428	 => "01001110001000010000011000010111",
		429	 => "01001110010010001101000011011100",
		430	 => "01001110011100001000111110001111",
		431	 => "01001110100110000100001000101001",
		432	 => "01001110101111111110100010100100",
		433	 => "01001110111001111000001011111010",
		434	 => "01001111000011110001000100100110",
		435	 => "01001111001101101001001100100000",
		436	 => "01001111010111100000100011100011",
		437	 => "01001111100001010111001001101000",
		438	 => "01001111101011001100111110101010",
		439	 => "01001111110101000010000010100011",
		440	 => "01001111111110110110010101001101",
		441	 => "01010000001000101001110110100000",
		442	 => "01010000010010011100100110011000",
		443	 => "01010000011100001110100100101111",
		444	 => "01010000100101111111110001011110",
		445	 => "01010000101111110000001100011111",
		446	 => "01010000111001011111110101101100",
		447	 => "01010001000011001110101101000000",
		448	 => "01010001001100111100110010010100",
		449	 => "01010001010110101010000101100010",
		450	 => "01010001100000010110100110100100",
		451	 => "01010001101010000010010101010101",
		452	 => "01010001110011101101010001101110",
		453	 => "01010001111101010111011011101001",
		454	 => "01010010000111000000110011000001",
		455	 => "01010010010000101001010111101111",
		456	 => "01010010011010010001001001101110",
		457	 => "01010010100011111000001000110111",
		458	 => "01010010101101011110010101000101",
		459	 => "01010010110111000011101110010010",
		460	 => "01010011000000101000010100010111",
		461	 => "01010011001010001100000111010000",
		462	 => "01010011010011101111000110110101",
		463	 => "01010011011101010001010011000001",
		464	 => "01010011100110110010101011101111",
		465	 => "01010011110000010011010000111000",
		466	 => "01010011111001110011000010010111",
		467	 => "01010100000011010010000000000101",
		468	 => "01010100001100110000001001111101",
		469	 => "01010100010110001101011111111001",
		470	 => "01010100011111101010000001110011",
		471	 => "01010100101001000101101111100101",
		472	 => "01010100110010100000101001001010",
		473	 => "01010100111011111010101110011100",
		474	 => "01010101000101010011111111010100",
		475	 => "01010101001110101100011011101101",
		476	 => "01010101011000000100000011100010",
		477	 => "01010101100001011010110110101100",
		478	 => "01010101101010110000110101000110",
		479	 => "01010101110100000101111110101010",
		480	 => "01010101111101011010010011010010",
		481	 => "01010110000110101101110010111000",
		482	 => "01010110010000000000011101010111",
		483	 => "01010110011001010010010010101010",
		484	 => "01010110100010100011010010101001",
		485	 => "01010110101011110011011101010000",
		486	 => "01010110110101000010110010011001",
		487	 => "01010110111110010001010001111110",
		488	 => "01010111000111011110111011111001",
		489	 => "01010111010000101011110000000101",
		490	 => "01010111011001110111101110011100",
		491	 => "01010111100011000010110110111001",
		492	 => "01010111101100001101001001010110",
		493	 => "01010111110101010110100101101100",
		494	 => "01010111111110011111001011110111",
		495	 => "01011000000111100110111011110001",
		496	 => "01011000010000101101110101010100",
		497	 => "01011000011001110011111000011011",
		498	 => "01011000100010111001000100111111",
		499	 => "01011000101011111101011010111100",
		500	 => "01011000110101000000111010001100",
		501	 => "01011000111110000011100010101001",
		502	 => "01011001000111000101010100001101",
		503	 => "01011001010000000110001110110100",
		504	 => "01011001011001000110010010010111",
		505	 => "01011001100010000101011110110001",
		506	 => "01011001101011000011110011111101",
		507	 => "01011001110100000001010001110100",
		508	 => "01011001111100111101111000010010",
		509	 => "01011010000101111001100111010000",
		510	 => "01011010001110110100011110101010",
		511	 => "01011010010111101110011110011010",
		512	 => "01011010100000100111100110011001",
		513	 => "01011010101001011111110110100100",
		514	 => "01011010110010010111001110110100",
		515	 => "01011010111011001101101111000100",
		516	 => "01011011000100000011010111001111",
		517	 => "01011011001100111000000111001110",
		518	 => "01011011010101101011111110111101",
		519	 => "01011011011110011110111110010110",
		520	 => "01011011100111010001000101010011",
		521	 => "01011011110000000010010011110000",
		522	 => "01011011111000110010101001100111",
		523	 => "01011100000001100010000110110010",
		524	 => "01011100001010010000101011001100",
		525	 => "01011100010010111110010110110000",
		526	 => "01011100011011101011001001011000",
		527	 => "01011100100100010111000010111111",
		528	 => "01011100101101000010000011011111",
		529	 => "01011100110101101100001010110100",
		530	 => "01011100111110010101011000111000",
		531	 => "01011101000110111101101101100101",
		532	 => "01011101001111100101001000110110",
		533	 => "01011101011000001011101010100110",
		534	 => "01011101100000110001010010110000",
		535	 => "01011101101001010110000001001110",
		536	 => "01011101110001111001110101111100",
		537	 => "01011101111010011100110000110010",
		538	 => "01011110000010111110110001101110",
		539	 => "01011110001011011111111000101000",
		540	 => "01011110010100000000000101011101",
		541	 => "01011110011100011111011000000110",
		542	 => "01011110100100111101110000011110",
		543	 => "01011110101101011011001110100001",
		544	 => "01011110110101110111110010001001",
		545	 => "01011110111110010011011011010001",
		546	 => "01011111000110101110001001110011",
		547	 => "01011111001111000111111101101011",
		548	 => "01011111010111100000110110110011",
		549	 => "01011111011111111000110101000101",
		550	 => "01011111101000001111111000011110",
		551	 => "01011111110000100110000000111000",
		552	 => "01011111111000111011001110001101",
		553	 => "01100000000001001111100000011000",
		554	 => "01100000001001100010110111010101",
		555	 => "01100000010001110101010010111110",
		556	 => "01100000011010000110110011001110",
		557	 => "01100000100010010111011000000000",
		558	 => "01100000101010100111000001001111",
		559	 => "01100000110010110101101110110110",
		560	 => "01100000111011000011100000101111",
		561	 => "01100001000011010000010110110111",
		562	 => "01100001001011011100010001000110",
		563	 => "01100001010011100111001111011001",
		564	 => "01100001011011110001010001101011",
		565	 => "01100001100011111010010111110110",
		566	 => "01100001101100000010100001110110",
		567	 => "01100001110100001001101111100101",
		568	 => "01100001111100010000000000111110",
		569	 => "01100010000100010101010101111101",
		570	 => "01100010001100011001101110011101",
		571	 => "01100010010100011101001010010111",
		572	 => "01100010011100011111101001101001",
		573	 => "01100010100100100001001100001100",
		574	 => "01100010101100100001110001111011",
		575	 => "01100010110100100001011010110010",
		576	 => "01100010111100100000000110101100",
		577	 => "01100011000100011101110101100011",
		578	 => "01100011001100011010100111010100",
		579	 => "01100011010100010110011011111000",
		580	 => "01100011011100010001010011001100",
		581	 => "01100011100100001011001101001010",
		582	 => "01100011101100000100001001101101",
		583	 => "01100011110011111100001000110000",
		584	 => "01100011111011110011001010001111",
		585	 => "01100100000011101001001110000101",
		586	 => "01100100001011011110010100001101",
		587	 => "01100100010011010010011100100010",
		588	 => "01100100011011000101100110111111",
		589	 => "01100100100010110111110011011111",
		590	 => "01100100101010101001000001111111",
		591	 => "01100100110010011001010010011000",
		592	 => "01100100111010001000100100100110",
		593	 => "01100101000001110110111000100100",
		594	 => "01100101001001100100001110001110",
		595	 => "01100101010001010000100101011111",
		596	 => "01100101011000111011111110010010",
		597	 => "01100101100000100110011000100010",
		598	 => "01100101101000001111110100001010",
		599	 => "01100101101111111000010001000111",
		600	 => "01100101110111011111101111010011",
		601	 => "01100101111111000110001110101001",
		602	 => "01100110000110101011101111000101",
		603	 => "01100110001110010000010000100010",
		604	 => "01100110010101110011110010111011",
		605	 => "01100110011101010110010110001100",
		606	 => "01100110100100110111111010010000",
		607	 => "01100110101100011000011111000011",
		608	 => "01100110110011111000000100011111",
		609	 => "01100110111011010110101010100001",
		610	 => "01100111000010110100010001000011",
		611	 => "01100111001010010000111000000010",
		612	 => "01100111010001101100011111010111",
		613	 => "01100111011001000111000111000000",
		614	 => "01100111100000100000101110110110",
		615	 => "01100111100111111001010110110111",
		616	 => "01100111101111010000111110111100",
		617	 => "01100111110110100111100111000010",
		618	 => "01100111111101111101001111000100",
		619	 => "01101000000101010001110110111110",
		620	 => "01101000001100100101011110101010",
		621	 => "01101000010011111000000110000101",
		622	 => "01101000011011001001101101001011",
		623	 => "01101000100010011010010011110101",
		624	 => "01101000101001101001111010000001",
		625	 => "01101000110000111000011111101001",
		626	 => "01101000111000000110000100101001",
		627	 => "01101000111111010010101000111101",
		628	 => "01101001000110011110001100100000",
		629	 => "01101001001101101000101111001110",
		630	 => "01101001010100110010010001000010",
		631	 => "01101001011011111010110001111000",
		632	 => "01101001100011000010010001101100",
		633	 => "01101001101010001000110000011000",
		634	 => "01101001110001001110001101111010",
		635	 => "01101001111000010010101010001100",
		636	 => "01101001111111010110000101001010",
		637	 => "01101010000110011000011110110000",
		638	 => "01101010001101011001110110111001",
		639	 => "01101010010100011010001101100001",
		640	 => "01101010011011011001100010100100",
		641	 => "01101010100010010111110101111101",
		642	 => "01101010101001010101000111101000",
		643	 => "01101010110000010001010111100001",
		644	 => "01101010110111001100100101100100",
		645	 => "01101010111110000110110001101100",
		646	 => "01101011000100111111111011110100",
		647	 => "01101011001011111000000011111010",
		648	 => "01101011010010101111001001111000",
		649	 => "01101011011001100101001101101010",
		650	 => "01101011100000011010001111001101",
		651	 => "01101011100111001110001110011011",
		652	 => "01101011101110000001001011010000",
		653	 => "01101011110100110011000101101010",
		654	 => "01101011111011100011111101100010",
		655	 => "01101100000010010011110010110101",
		656	 => "01101100001001000010100101100000",
		657	 => "01101100001111110000010101011101",
		658	 => "01101100010110011101000010101001",
		659	 => "01101100011101001000101100111111",
		660	 => "01101100100011110011010100011100",
		661	 => "01101100101010011100111000111010",
		662	 => "01101100110001000101011010010111",
		663	 => "01101100110111101100111000101110",
		664	 => "01101100111110010011010011111011",
		665	 => "01101101000100111000101011111010",
		666	 => "01101101001011011101000000100111",
		667	 => "01101101010010000000010001111110",
		668	 => "01101101011000100010011111111010",
		669	 => "01101101011111000011101010011000",
		670	 => "01101101100101100011110001010011",
		671	 => "01101101101100000010110100101001",
		672	 => "01101101110010100000110100010100",
		673	 => "01101101111000111101110000010001",
		674	 => "01101101111111011001101000011011",
		675	 => "01101110000101110100011100101111",
		676	 => "01101110001100001110001101001001",
		677	 => "01101110010010100110111001100101",
		678	 => "01101110011000111110100001111111",
		679	 => "01101110011111010101000110010011",
		680	 => "01101110100101101010100110011100",
		681	 => "01101110101011111111000010011000",
		682	 => "01101110110010010010011010000010",
		683	 => "01101110111000100100101101010111",
		684	 => "01101110111110110101111100010010",
		685	 => "01101111000101000110000110101111",
		686	 => "01101111001011010101001100101100",
		687	 => "01101111010001100011001110000011",
		688	 => "01101111010111110000001010110001",
		689	 => "01101111011101111100000010110011",
		690	 => "01101111100100000110110110000100",
		691	 => "01101111101010010000100100100000",
		692	 => "01101111110000011001001110000101",
		693	 => "01101111110110100000110010101101",
		694	 => "01101111111100100111010010010110",
		695	 => "01110000000010101100101100111011",
		696	 => "01110000001000110001000010011001",
		697	 => "01110000001110110100010010101100",
		698	 => "01110000010100110110011101110001",
		699	 => "01110000011010110111100011100010",
		700	 => "01110000100000110111100011111110",
		701	 => "01110000100110110110011111000000",
		702	 => "01110000101100110100010100100100",
		703	 => "01110000110010110001000100100111",
		704	 => "01110000111000101100101111000110",
		705	 => "01110000111110100111010011111011",
		706	 => "01110001000100100000110011000101",
		707	 => "01110001001010011001001100011110",
		708	 => "01110001010000010000100000000100",
		709	 => "01110001010110000110101101110011",
		710	 => "01110001011011111011110101100111",
		711	 => "01110001100001101111110111011101",
		712	 => "01110001100111100010110011010010",
		713	 => "01110001101101010100101001000000",
		714	 => "01110001110011000101011000100110",
		715	 => "01110001111000110101000001111111",
		716	 => "01110001111110100011100101001000",
		717	 => "01110010000100010001000001111101",
		718	 => "01110010001001111101011000011100",
		719	 => "01110010001111101000101000011111",
		720	 => "01110010010101010010110010000100",
		721	 => "01110010011010111011110101001000",
		722	 => "01110010100000100011110001100110",
		723	 => "01110010100110001010100111011100",
		724	 => "01110010101011110000010110100110",
		725	 => "01110010110001010100111111000000",
		726	 => "01110010110110111000100000101000",
		727	 => "01110010111100011010111011011000",
		728	 => "01110011000001111100001111001111",
		729	 => "01110011000111011100011100001001",
		730	 => "01110011001100111011100010000011",
		731	 => "01110011010010011001100000111000",
		732	 => "01110011010111110110011000100110",
		733	 => "01110011011101010010001001001001",
		734	 => "01110011100010101100110010011110",
		735	 => "01110011101000000110010100100010",
		736	 => "01110011101101011110101111010000",
		737	 => "01110011110010110110000010100111",
		738	 => "01110011111000001100001110100011",
		739	 => "01110011111101100001010010111111",
		740	 => "01110100000010110101001111111010",
		741	 => "01110100001000001000000101010000",
		742	 => "01110100001101011001110010111101",
		743	 => "01110100010010101010011000111110",
		744	 => "01110100010111111001110111010000",
		745	 => "01110100011101001000001101110001",
		746	 => "01110100100010010101011100011011",
		747	 => "01110100100111100001100011001101",
		748	 => "01110100101100101100100010000011",
		749	 => "01110100110001110110011000111010",
		750	 => "01110100110110111111000111101111",
		751	 => "01110100111100000110101110011110",
		752	 => "01110101000001001101001101000101",
		753	 => "01110101000110010010100011100000",
		754	 => "01110101001011010110110001101100",
		755	 => "01110101010000011001110111100110",
		756	 => "01110101010101011011110101001011",
		757	 => "01110101011010011100101010011000",
		758	 => "01110101011111011100010111001010",
		759	 => "01110101100100011010111011011101",
		760	 => "01110101101001011000010111001111",
		761	 => "01110101101110010100101010011100",
		762	 => "01110101110011001111110101000010",
		763	 => "01110101111000001001110110111101",
		764	 => "01110101111101000010110000001010",
		765	 => "01110110000001111010100000100111",
		766	 => "01110110000110110001001000010001",
		767	 => "01110110001011100110100111000011",
		768	 => "01110110010000011010111100111100",
		769	 => "01110110010101001110001001111001",
		770	 => "01110110011010000000001101110110",
		771	 => "01110110011110110001001000110000",
		772	 => "01110110100011100000111010100101",
		773	 => "01110110101000001111100011010010",
		774	 => "01110110101100111101000010110011",
		775	 => "01110110110001101001011001000110",
		776	 => "01110110110110010100100110001000",
		777	 => "01110110111010111110101001110111",
		778	 => "01110110111111100111100100001110",
		779	 => "01110111000100001111010101001011",
		780	 => "01110111001000110101111100101101",
		781	 => "01110111001101011011011010101110",
		782	 => "01110111010001111111101111001110",
		783	 => "01110111010110100010111010001000",
		784	 => "01110111011011000100111011011011",
		785	 => "01110111011111100101110011000011",
		786	 => "01110111100100000101100000111101",
		787	 => "01110111101000100100000101001000",
		788	 => "01110111101101000001011111011111",
		789	 => "01110111110001011101110000000001",
		790	 => "01110111110101111000110110101010",
		791	 => "01110111111010010010110011011000",
		792	 => "01110111111110101011100110001000",
		793	 => "01111000000011000011001110111000",
		794	 => "01111000000111011001101101100100",
		795	 => "01111000001011101111000010001010",
		796	 => "01111000010000000011001100101000",
		797	 => "01111000010100010110001100111011",
		798	 => "01111000011000101000000010111111",
		799	 => "01111000011100111000101110110011",
		800	 => "01111000100001001000010000010011",
		801	 => "01111000100101010110100111011110",
		802	 => "01111000101001100011110100010000",
		803	 => "01111000101101101111110110101000",
		804	 => "01111000110001111010101110100001",
		805	 => "01111000110110000100011011111011",
		806	 => "01111000111010001100111110110001",
		807	 => "01111000111110010100010111000011",
		808	 => "01111001000010011010100100101100",
		809	 => "01111001000110011111100111101011",
		810	 => "01111001001010100011011111111110",
		811	 => "01111001001110100110001101100000",
		812	 => "01111001010010100111110000010001",
		813	 => "01111001010110101000001000001110",
		814	 => "01111001011010100111010101010100",
		815	 => "01111001011110100101010111100000",
		816	 => "01111001100010100010001110110001",
		817	 => "01111001100110011101111011000011",
		818	 => "01111001101010011000011100010101",
		819	 => "01111001101110010001110010100100",
		820	 => "01111001110010001001111101101101",
		821	 => "01111001110110000000111101101111",
		822	 => "01111001111001110110110010100110",
		823	 => "01111001111101101011011100010001",
		824	 => "01111010000001011110111010101101",
		825	 => "01111010000101010001001101110111",
		826	 => "01111010001001000010010101101110",
		827	 => "01111010001100110010010010001111",
		828	 => "01111010010000100001000011011000",
		829	 => "01111010010100001110101001000110",
		830	 => "01111010010111111011000011011000",
		831	 => "01111010011011100110010010001010",
		832	 => "01111010011111010000010101011011",
		833	 => "01111010100010111001001101001000",
		834	 => "01111010100110100000111001001111",
		835	 => "01111010101010000111011001101110",
		836	 => "01111010101101101100101110100011",
		837	 => "01111010110001010000110111101011",
		838	 => "01111010110100110011110101000101",
		839	 => "01111010111000010101100110101110",
		840	 => "01111010111011110110001100100011",
		841	 => "01111010111111010101100110100011",
		842	 => "01111011000010110011110100101100",
		843	 => "01111011000110010000110110111011",
		844	 => "01111011001001101100101101001111",
		845	 => "01111011001101000111010111100100",
		846	 => "01111011010000100000110101111010",
		847	 => "01111011010011111001001000001110",
		848	 => "01111011010111010000001110011101",
		849	 => "01111011011010100110001000100110",
		850	 => "01111011011101111010110110101000",
		851	 => "01111011100001001110011000011110",
		852	 => "01111011100100100000101110001001",
		853	 => "01111011100111110001110111100101",
		854	 => "01111011101011000001110100110001",
		855	 => "01111011101110010000100101101010",
		856	 => "01111011110001011110001010001111",
		857	 => "01111011110100101010100010011110",
		858	 => "01111011110111110101101110010100",
		859	 => "01111011111010111111101101110000",
		860	 => "01111011111110001000100000110000",
		861	 => "01111100000001010000000111010001",
		862	 => "01111100000100010110100001010011",
		863	 => "01111100000111011011101110110010",
		864	 => "01111100001010011111101111101110",
		865	 => "01111100001101100010100100000100",
		866	 => "01111100010000100100001011110010",
		867	 => "01111100010011100100100110110110",
		868	 => "01111100010110100011110101001111",
		869	 => "01111100011001100001110110111011",
		870	 => "01111100011100011110101011111000",
		871	 => "01111100011111011010010100000100",
		872	 => "01111100100010010100101111011101",
		873	 => "01111100100101001101111110000010",
		874	 => "01111100101000000101111111110001",
		875	 => "01111100101010111100110100100111",
		876	 => "01111100101101110010011100100100",
		877	 => "01111100110000100110110111100101",
		878	 => "01111100110011011010000101101000",
		879	 => "01111100110110001100000110101101",
		880	 => "01111100111000111100111010110001",
		881	 => "01111100111011101100100001110011",
		882	 => "01111100111110011010111011110000",
		883	 => "01111101000001001000001000100111",
		884	 => "01111101000011110100001000010111",
		885	 => "01111101000110011110111010111110",
		886	 => "01111101001001001000100000011010",
		887	 => "01111101001011110000111000101010",
		888	 => "01111101001110011000000011101100",
		889	 => "01111101010000111110000001011110",
		890	 => "01111101010011100010110001111110",
		891	 => "01111101010110000110010101001100",
		892	 => "01111101011000101000101011000101",
		893	 => "01111101011011001001110011101001",
		894	 => "01111101011101101001101110110101",
		895	 => "01111101100000001000011100100111",
		896	 => "01111101100010100101111100111111",
		897	 => "01111101100101000010001111111011",
		898	 => "01111101100111011101010101011010",
		899	 => "01111101101001110111001101011001",
		900	 => "01111101101100001111110111110111",
		901	 => "01111101101110100111010100110100",
		902	 => "01111101110000111101100100001101",
		903	 => "01111101110011010010100110000001",
		904	 => "01111101110101100110011010001110",
		905	 => "01111101110111111001000000110100",
		906	 => "01111101111010001010011001110000",
		907	 => "01111101111100011010100101000010",
		908	 => "01111101111110101001100010100111",
		909	 => "01111110000000110111010010011111",
		910	 => "01111110000011000011110100101001",
		911	 => "01111110000101001111001001000010",
		912	 => "01111110000111011001001111101001",
		913	 => "01111110001001100010001000011110",
		914	 => "01111110001011101001110011011111",
		915	 => "01111110001101110000010000101010",
		916	 => "01111110001111110101011111111110",
		917	 => "01111110010001111001100001011011",
		918	 => "01111110010011111100010100111110",
		919	 => "01111110010101111101111010100110",
		920	 => "01111110010111111110010010010011",
		921	 => "01111110011001111101011100000010",
		922	 => "01111110011011111011010111110011",
		923	 => "01111110011101111000000101100101",
		924	 => "01111110011111110011100101010110",
		925	 => "01111110100001101101110111000101",
		926	 => "01111110100011100110111010110001",
		927	 => "01111110100101011110110000011001",
		928	 => "01111110100111010101010111111100",
		929	 => "01111110101001001010110001011000",
		930	 => "01111110101010111110111100101100",
		931	 => "01111110101100110001111001110111",
		932	 => "01111110101110100011101000111001",
		933	 => "01111110110000010100001001101111",
		934	 => "01111110110010000011011100011010",
		935	 => "01111110110011110001100000110111",
		936	 => "01111110110101011110010111000110",
		937	 => "01111110110111001001111111000110",
		938	 => "01111110111000110100011000110101",
		939	 => "01111110111010011101100100010011",
		940	 => "01111110111100000101100001011111",
		941	 => "01111110111101101100010000011000",
		942	 => "01111110111111010001110000111100",
		943	 => "01111111000000110110000011001010",
		944	 => "01111111000010011001000111000011",
		945	 => "01111111000011111010111100100100",
		946	 => "01111111000101011011100011101101",
		947	 => "01111111000110111010111100011101",
		948	 => "01111111001000011001000110110011",
		949	 => "01111111001001110110000010101111",
		950	 => "01111111001011010001110000001110",
		951	 => "01111111001100101100001111010000",
		952	 => "01111111001110000101011111110101",
		953	 => "01111111001111011101100001111100",
		954	 => "01111111010000110100010101100011",
		955	 => "01111111010010001001111010101010",
		956	 => "01111111010011011110010001010000",
		957	 => "01111111010100110001011001010100",
		958	 => "01111111010110000011010010110110",
		959	 => "01111111010111010011111101110101",
		960	 => "01111111011000100011011010001111",
		961	 => "01111111011001110001101000000100",
		962	 => "01111111011010111110100111010100",
		963	 => "01111111011100001010010111111101",
		964	 => "01111111011101010100111001111111",
		965	 => "01111111011110011110001101011010",
		966	 => "01111111011111100110010010001011",
		967	 => "01111111100000101101001000010100",
		968	 => "01111111100001110010101111110010",
		969	 => "01111111100010110111001000100110",
		970	 => "01111111100011111010010010101111",
		971	 => "01111111100100111100001110001100",
		972	 => "01111111100101111100111010111100",
		973	 => "01111111100110111100011000111111",
		974	 => "01111111100111111010101000010101",
		975	 => "01111111101000110111101000111100",
		976	 => "01111111101001110011011010110100",
		977	 => "01111111101010101101111101111100",
		978	 => "01111111101011100111010010010100",
		979	 => "01111111101100011111010111111100",
		980	 => "01111111101101010110001110110010",
		981	 => "01111111101110001011110110110111",
		982	 => "01111111101111000000010000001010",
		983	 => "01111111101111110011011010101001",
		984	 => "01111111110000100101010110010110",
		985	 => "01111111110001010110000011001110",
		986	 => "01111111110010000101100001010011",
		987	 => "01111111110010110011110000100011",
		988	 => "01111111110011100000110000111110",
		989	 => "01111111110100001100100010100011",
		990	 => "01111111110100110111000101010010",
		991	 => "01111111110101100000011001001011",
		992	 => "01111111110110001000011110001101",
		993	 => "01111111110110101111010100011000",
		994	 => "01111111110111010100111011101100",
		995	 => "01111111110111111001010100001000",
		996	 => "01111111111000011100011101101011",
		997	 => "01111111111000111110011000010110",
		998	 => "01111111111001011111000100001000",
		999	 => "01111111111001111110100001000000",
		1000	 => "01111111111010011100101110111111",
		1001	 => "01111111111010111001101110000101",
		1002	 => "01111111111011010101011110010000",
		1003	 => "01111111111011101111111111100001",
		1004	 => "01111111111100001001010001110111",
		1005	 => "01111111111100100001010101010011",
		1006	 => "01111111111100111000001001110011",
		1007	 => "01111111111101001101101111011000",
		1008	 => "01111111111101100010000110000010",
		1009	 => "01111111111101110101001101101111",
		1010	 => "01111111111110000111000110100001",
		1011	 => "01111111111110010111110000010111",
		1012	 => "01111111111110100111001011010001",
		1013	 => "01111111111110110101010111001110",
		1014	 => "01111111111111000010010100001111",
		1015	 => "01111111111111001110000010010011",
		1016	 => "01111111111111011000100001011010",
		1017	 => "01111111111111100001110001100100",
		1018	 => "01111111111111101001110010110010",
		1019	 => "01111111111111110000100101000010",
		1020	 => "01111111111111110110001000010110",
		1021	 => "01111111111111111010011100101100",
		1022	 => "01111111111111111101100010000101",
		1023	 => "01111111111111111111011000100001");

end wave_rom_package;

